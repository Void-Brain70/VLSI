module main;

initial 

begin

$display("anik das");

$finish ;

end

endmodule